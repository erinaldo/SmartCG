<?xml version="1.0" standalone="yes"?>
<Formulario>
  <Cabecera>
    <Codigo>MISIIDATL</Codigo>
    <Descripcion>demo consulta local 1</Descripcion>
  </Cabecera>
  <Control>
    <Nombre>cmbClaveOperacion</Nombre>
    <Tipo>ComboBox</Tipo>
    <Valor />
  </Control>
  <Control>
    <Nombre>txtMaskFechaExpedicion</Nombre>
    <Tipo>MaskedTextBox</Tipo>
    <Valor />
  </Control>
  <Control>
    <Nombre>rbEstadoPdteEnvio</Nombre>
    <Tipo>RadioButton</Tipo>
    <Valor>0</Valor>
  </Control>
  <Control>
    <Nombre>rbEstadoAceptadoErrores</Nombre>
    <Tipo>RadioButton</Tipo>
    <Valor>0</Valor>
  </Control>
  <Control>
    <Nombre>rbEstadoCorrecto</Nombre>
    <Tipo>RadioButton</Tipo>
    <Valor>0</Valor>
  </Control>
  <Control>
    <Nombre>rbEstadoSoloErrores</Nombre>
    <Tipo>RadioButton</Tipo>
    <Valor>0</Valor>
  </Control>
  <Control>
    <Nombre>rbEstadoTodas</Nombre>
    <Tipo>RadioButton</Tipo>
    <Valor>1</Valor>
  </Control>
  <Control>
    <Nombre>txtNumSerieFactura</Nombre>
    <Tipo>TextBox</Tipo>
    <Valor />
  </Control>
  <Control>
    <Nombre>cmbTipoIdentif</Nombre>
    <Tipo>ComboBox</Tipo>
    <Valor />
  </Control>
  <Control>
    <Nombre>txtNombreRazon</Nombre>
    <Tipo>TextBox</Tipo>
    <Valor />
  </Control>
  <Control>
    <Nombre>txtCodPais</Nombre>
    <Tipo>TextBox</Tipo>
    <Valor />
  </Control>
  <Control>
    <Nombre>txtNIF</Nombre>
    <Tipo>TextBox</Tipo>
    <Valor />
  </Control>
  <Control>
    <Nombre>rbOtro</Nombre>
    <Tipo>RadioButton</Tipo>
    <Valor>0</Valor>
  </Control>
  <Control>
    <Nombre>rbNIF</Nombre>
    <Tipo>RadioButton</Tipo>
    <Valor>1</Valor>
  </Control>
  <Control>
    <Nombre>txtEjercicio</Nombre>
    <Tipo>TextBox</Tipo>
    <Valor>2017</Valor>
  </Control>
  <Control>
    <Nombre>tgTexBoxSelCiaFiscal</Nombre>
    <Tipo>TGTexBoxSel</Tipo>
    <Valor>SA - CONTA, S.L. - B61350765</Valor>
  </Control>
  <Control>
    <Nombre>txtElemento</Nombre>
    <Tipo>TextBox</Tipo>
    <Valor>SA - CONTA, S.L. - B61350765</Valor>
  </Control>
  <Control>
    <Nombre>cmbPeriodo</Nombre>
    <Tipo>ComboBox</Tipo>
    <Valor>04</Valor>
  </Control>
  <Control>
    <Nombre>cmbLibro</Nombre>
    <Tipo>ComboBox</Tipo>
    <Valor>03</Valor>
  </Control>
  <Control>
    <Nombre>txtLibroDesc</Nombre>
    <Tipo>TextBox</Tipo>
    <Valor>Facturas Recibidas</Valor>
  </Control>
</Formulario>